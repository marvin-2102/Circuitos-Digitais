IBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SAIDABC IS

	PORT(CK, RST, WR, RD, EM, FU: IN STD_LOGIC;
		  EN_R, EN_W: OUT STD_LOGIC;
		  Q: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	    );


END SAIDABC;


ARCHITECTURE MOORE OF SAIDABC IS
	
	
COMPONENT MDE 	

	PORT(CK, RST, WR, RD, EM, FU: IN STD_LOGIC;
		  Q: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	    );

END COMPONENT;

SIGNAL S: STD_lOGIC_VECTOR(1 DOWNTO 0);

BEGIN

M0: MDE PORT MAP(CK, RST, WR, RD, EM, FU, S);


Q <= S;
EN_W <= NOT S(0) AND S(1);
EN_R <= S(0) AND NOT S(1);


END MOORE;