LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MDE IS

	PORT(CK, RST, WR, RD, EM, FU: IN STD_LOGIC;
		  Q: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	    );


END MDE;


ARCHITECTURE MOORE OF MDE IS
	TYPE ST IS (ESPERAR, LER, ESCREVER);
	SIGNAL ESTADO: ST;

BEGIN
	PROCESS(CK, RST)
	BEGIN
		IF(RST = '1' AND RD = '0' AND WR = '0') THEN
			ESTADO <= ESPERAR;
		ELSIF(CK'EVENT AND CK = '1') THEN
			CASE ESTADO IS
				WHEN ESPERAR =>
					IF(WR = '1' AND RD = '0' AND FU = '0') THEN ESTADO <= ESCREVER;
					ELSIF(WR = '0' AND RD = '1' AND EM = '0') THEN ESTADO <= LER;
						END IF;
				WHEN LER =>
					IF CK = '1' THEN ESTADO <= ESPERAR;
					END IF;
				WHEN ESCREVER =>
					IF CK = '1' THEN ESTADO <= ESPERAR; 
					END IF;
			END CASE;
		END IF;
	END PROCESS;
	
	WITH ESTADO SELECT
		Q <= "00" WHEN ESPERAR, 
		     "01" WHEN LER,
			  "10" WHEN ESCREVER;
END MOORE;
